// decodes 10b symbols into the 8b control/data character
// takes data in the order abcdei fghj
// input_data -> output_data is a combinational path

module decoder_8b10b (
  input  logic [9:0] input_data,
  output logic [7:0] output_data,
  output logic [7:0] output_ctrl
);
  logic [9:0] rom_addr;
  logic [8:0] krom_read;
  logic [8:0] drom_read;

  logic [8:0] krom [1023:0];
  logic [8:0] drom [1023:0];

  assign rom_addr = input_data;
  assign krom_read = krom[rom_addr];
  assign drom_read = drom[rom_addr];
  assign output_data = drom_read[7:0];
  assign output_ctrl = krom_read[7:0];
  
  initial begin
    krom[85] = 9'b110110111;
    krom[86] = 9'b100110111;
    krom[87] = 9'b111110111;
    krom[89] = 9'b111010111;
    krom[90] = 9'b101010111;
    krom[91] = 9'b100010111;
    krom[92] = 9'b101110111;
    krom[93] = 9'b110010111;
    krom[101] = 9'b110101000;
    krom[102] = 9'b100101000;
    krom[103] = 9'b111101000;
    krom[105] = 9'b111001000;
    krom[106] = 9'b101001000;
    krom[107] = 9'b100001000;
    krom[108] = 9'b101101000;
    krom[109] = 9'b110001000;
    krom[114] = 9'b110000111;
    krom[115] = 9'b101100111;
    krom[116] = 9'b100000111;
    krom[117] = 9'b101000111;
    krom[118] = 9'b111000111;
    krom[120] = 9'b111100111;
    krom[121] = 9'b100100111;
    krom[122] = 9'b110100111;
    krom[149] = 9'b110111011;
    krom[150] = 9'b100111011;
    krom[151] = 9'b111111011;
    krom[153] = 9'b111011011;
    krom[154] = 9'b101011011;
    krom[155] = 9'b100011011;
    krom[156] = 9'b101111011;
    krom[157] = 9'b110011011;
    krom[165] = 9'b110100100;
    krom[166] = 9'b100100100;
    krom[167] = 9'b111100100;
    krom[169] = 9'b111000100;
    krom[170] = 9'b101000100;
    krom[171] = 9'b100000100;
    krom[172] = 9'b101100100;
    krom[173] = 9'b110000100;
    krom[178] = 9'b110010100;
    krom[179] = 9'b101110100;
    krom[180] = 9'b100010100;
    krom[181] = 9'b101010100;
    krom[182] = 9'b111010100;
    krom[183] = 9'b011110100;
    krom[184] = 9'b111110100;
    krom[185] = 9'b100110100;
    krom[186] = 9'b110110100;
    krom[187] = 9'b000010100;
    krom[188] = 9'b001110100;
    krom[189] = 9'b010010100;
    krom[197] = 9'b110111000;
    krom[198] = 9'b100111000;
    krom[199] = 9'b111111000;
    krom[201] = 9'b111011000;
    krom[202] = 9'b101011000;
    krom[203] = 9'b100011000;
    krom[204] = 9'b101111000;
    krom[205] = 9'b110011000;
    krom[210] = 9'b110001100;
    krom[211] = 9'b101101100;
    krom[212] = 9'b100001100;
    krom[213] = 9'b101001100;
    krom[214] = 9'b111001100;
    krom[215] = 9'b011101100;
    krom[216] = 9'b111101100;
    krom[217] = 9'b100101100;
    krom[218] = 9'b110101100;
    krom[219] = 9'b000001100;
    krom[220] = 9'b001101100;
    krom[221] = 9'b010001100;
    krom[242] = 9'b010011100;
    krom[243] = 9'b001111100;
    krom[244] = 9'b000011100;
    krom[245] = 9'b001011100;
    krom[246] = 9'b011011100;
    krom[248] = 9'b011111100;
    krom[249] = 9'b000111100;
    krom[250] = 9'b010111100;
    krom[277] = 9'b110111101;
    krom[278] = 9'b100111101;
    krom[279] = 9'b111111101;
    krom[281] = 9'b111011101;
    krom[282] = 9'b101011101;
    krom[283] = 9'b100011101;
    krom[284] = 9'b101111101;
    krom[285] = 9'b110011101;
    krom[293] = 9'b110100010;
    krom[294] = 9'b100100010;
    krom[295] = 9'b111100010;
    krom[297] = 9'b111000010;
    krom[298] = 9'b101000010;
    krom[299] = 9'b100000010;
    krom[300] = 9'b101100010;
    krom[301] = 9'b110000010;
    krom[306] = 9'b110010010;
    krom[307] = 9'b101110010;
    krom[308] = 9'b100010010;
    krom[309] = 9'b101010010;
    krom[310] = 9'b111010010;
    krom[311] = 9'b011110010;
    krom[312] = 9'b111110010;
    krom[313] = 9'b100110010;
    krom[314] = 9'b110110010;
    krom[315] = 9'b000010010;
    krom[316] = 9'b001110010;
    krom[317] = 9'b010010010;
    krom[325] = 9'b110111111;
    krom[326] = 9'b100111111;
    krom[327] = 9'b111111111;
    krom[329] = 9'b111011111;
    krom[330] = 9'b101011111;
    krom[331] = 9'b100011111;
    krom[332] = 9'b101111111;
    krom[333] = 9'b110011111;
    krom[338] = 9'b110001010;
    krom[339] = 9'b101101010;
    krom[340] = 9'b100001010;
    krom[341] = 9'b101001010;
    krom[342] = 9'b111001010;
    krom[343] = 9'b011101010;
    krom[344] = 9'b111101010;
    krom[345] = 9'b100101010;
    krom[346] = 9'b110101010;
    krom[347] = 9'b000001010;
    krom[348] = 9'b001101010;
    krom[349] = 9'b010001010;
    krom[354] = 9'b110011010;
    krom[355] = 9'b101111010;
    krom[356] = 9'b100011010;
    krom[357] = 9'b101011010;
    krom[358] = 9'b111011010;
    krom[359] = 9'b011111010;
    krom[360] = 9'b111111010;
    krom[361] = 9'b100111010;
    krom[362] = 9'b110111010;
    krom[363] = 9'b000011010;
    krom[364] = 9'b001111010;
    krom[365] = 9'b010011010;
    krom[370] = 9'b010001111;
    krom[371] = 9'b001101111;
    krom[372] = 9'b000001111;
    krom[373] = 9'b001001111;
    krom[374] = 9'b011001111;
    krom[376] = 9'b011101111;
    krom[377] = 9'b000101111;
    krom[378] = 9'b010101111;
    krom[389] = 9'b110100000;
    krom[390] = 9'b100100000;
    krom[391] = 9'b111100000;
    krom[393] = 9'b111000000;
    krom[394] = 9'b101000000;
    krom[395] = 9'b100000000;
    krom[396] = 9'b101100000;
    krom[397] = 9'b110000000;
    krom[402] = 9'b110000110;
    krom[403] = 9'b101100110;
    krom[404] = 9'b100000110;
    krom[405] = 9'b101000110;
    krom[406] = 9'b111000110;
    krom[407] = 9'b011100110;
    krom[408] = 9'b111100110;
    krom[409] = 9'b100100110;
    krom[410] = 9'b110100110;
    krom[411] = 9'b000000110;
    krom[412] = 9'b001100110;
    krom[413] = 9'b010000110;
    krom[418] = 9'b110010110;
    krom[419] = 9'b101110110;
    krom[420] = 9'b100010110;
    krom[421] = 9'b101010110;
    krom[422] = 9'b111010110;
    krom[423] = 9'b011110110;
    krom[424] = 9'b111110110;
    krom[425] = 9'b100110110;
    krom[426] = 9'b110110110;
    krom[427] = 9'b000010110;
    krom[428] = 9'b001110110;
    krom[429] = 9'b010010110;
    krom[434] = 9'b010010000;
    krom[435] = 9'b001110000;
    krom[436] = 9'b000010000;
    krom[437] = 9'b001010000;
    krom[438] = 9'b011010000;
    krom[440] = 9'b011110000;
    krom[441] = 9'b000110000;
    krom[442] = 9'b010110000;
    krom[450] = 9'b110001110;
    krom[451] = 9'b101101110;
    krom[452] = 9'b100001110;
    krom[453] = 9'b101001110;
    krom[454] = 9'b111001110;
    krom[455] = 9'b011101110;
    krom[456] = 9'b111101110;
    krom[457] = 9'b100101110;
    krom[458] = 9'b110101110;
    krom[459] = 9'b000001110;
    krom[460] = 9'b001101110;
    krom[461] = 9'b010001110;
    krom[466] = 9'b010000001;
    krom[467] = 9'b001100001;
    krom[468] = 9'b000000001;
    krom[469] = 9'b001000001;
    krom[470] = 9'b011000001;
    krom[472] = 9'b011100001;
    krom[473] = 9'b000100001;
    krom[474] = 9'b010100001;
    krom[482] = 9'b010011110;
    krom[483] = 9'b001111110;
    krom[484] = 9'b000011110;
    krom[485] = 9'b001011110;
    krom[486] = 9'b011011110;
    krom[488] = 9'b011111110;
    krom[489] = 9'b000111110;
    krom[490] = 9'b010111110;
    krom[533] = 9'b110111110;
    krom[534] = 9'b100111110;
    krom[535] = 9'b111111110;
    krom[537] = 9'b111011110;
    krom[538] = 9'b101011110;
    krom[539] = 9'b100011110;
    krom[540] = 9'b101111110;
    krom[541] = 9'b110011110;
    krom[549] = 9'b110100001;
    krom[550] = 9'b100100001;
    krom[551] = 9'b111100001;
    krom[553] = 9'b111000001;
    krom[554] = 9'b101000001;
    krom[555] = 9'b100000001;
    krom[556] = 9'b101100001;
    krom[557] = 9'b110000001;
    krom[562] = 9'b110010001;
    krom[563] = 9'b101110001;
    krom[564] = 9'b100010001;
    krom[565] = 9'b101010001;
    krom[566] = 9'b111010001;
    krom[567] = 9'b011110001;
    krom[568] = 9'b111110001;
    krom[569] = 9'b100110001;
    krom[570] = 9'b110110001;
    krom[571] = 9'b000010001;
    krom[572] = 9'b001110001;
    krom[573] = 9'b010010001;
    krom[581] = 9'b110110000;
    krom[582] = 9'b100110000;
    krom[583] = 9'b111110000;
    krom[585] = 9'b111010000;
    krom[586] = 9'b101010000;
    krom[587] = 9'b100010000;
    krom[588] = 9'b101110000;
    krom[589] = 9'b110010000;
    krom[594] = 9'b110001001;
    krom[595] = 9'b101101001;
    krom[596] = 9'b100001001;
    krom[597] = 9'b101001001;
    krom[598] = 9'b111001001;
    krom[599] = 9'b011101001;
    krom[600] = 9'b111101001;
    krom[601] = 9'b100101001;
    krom[602] = 9'b110101001;
    krom[603] = 9'b000001001;
    krom[604] = 9'b001101001;
    krom[605] = 9'b010001001;
    krom[610] = 9'b110011001;
    krom[611] = 9'b101111001;
    krom[612] = 9'b100011001;
    krom[613] = 9'b101011001;
    krom[614] = 9'b111011001;
    krom[615] = 9'b011111001;
    krom[616] = 9'b111111001;
    krom[617] = 9'b100111001;
    krom[618] = 9'b110111001;
    krom[619] = 9'b000011001;
    krom[620] = 9'b001111001;
    krom[621] = 9'b010011001;
    krom[626] = 9'b010000000;
    krom[627] = 9'b001100000;
    krom[628] = 9'b000000000;
    krom[629] = 9'b001000000;
    krom[630] = 9'b011000000;
    krom[632] = 9'b011100000;
    krom[633] = 9'b000100000;
    krom[634] = 9'b010100000;
    krom[645] = 9'b110101111;
    krom[646] = 9'b100101111;
    krom[647] = 9'b111101111;
    krom[649] = 9'b111001111;
    krom[650] = 9'b101001111;
    krom[651] = 9'b100001111;
    krom[652] = 9'b101101111;
    krom[653] = 9'b110001111;
    krom[658] = 9'b110000101;
    krom[659] = 9'b101100101;
    krom[660] = 9'b100000101;
    krom[661] = 9'b101000101;
    krom[662] = 9'b111000101;
    krom[663] = 9'b011100101;
    krom[664] = 9'b111100101;
    krom[665] = 9'b100100101;
    krom[666] = 9'b110100101;
    krom[667] = 9'b000000101;
    krom[668] = 9'b001100101;
    krom[669] = 9'b010000101;
    krom[674] = 9'b110010101;
    krom[675] = 9'b101110101;
    krom[676] = 9'b100010101;
    krom[677] = 9'b101010101;
    krom[678] = 9'b111010101;
    krom[679] = 9'b011110101;
    krom[680] = 9'b111110101;
    krom[681] = 9'b100110101;
    krom[682] = 9'b110110101;
    krom[683] = 9'b000010101;
    krom[684] = 9'b001110101;
    krom[685] = 9'b010010101;
    krom[690] = 9'b010011111;
    krom[691] = 9'b001111111;
    krom[692] = 9'b000011111;
    krom[693] = 9'b001011111;
    krom[694] = 9'b011011111;
    krom[696] = 9'b011111111;
    krom[697] = 9'b000111111;
    krom[698] = 9'b010111111;
    krom[706] = 9'b110001101;
    krom[707] = 9'b101101101;
    krom[708] = 9'b100001101;
    krom[709] = 9'b101001101;
    krom[710] = 9'b111001101;
    krom[711] = 9'b011101101;
    krom[712] = 9'b111101101;
    krom[713] = 9'b100101101;
    krom[714] = 9'b110101101;
    krom[715] = 9'b000001101;
    krom[716] = 9'b001101101;
    krom[717] = 9'b010001101;
    krom[722] = 9'b010000010;
    krom[723] = 9'b001100010;
    krom[724] = 9'b000000010;
    krom[725] = 9'b001000010;
    krom[726] = 9'b011000010;
    krom[728] = 9'b011100010;
    krom[729] = 9'b000100010;
    krom[730] = 9'b010100010;
    krom[738] = 9'b010011101;
    krom[739] = 9'b001111101;
    krom[740] = 9'b000011101;
    krom[741] = 9'b001011101;
    krom[742] = 9'b011011101;
    krom[744] = 9'b011111101;
    krom[745] = 9'b000111101;
    krom[746] = 9'b010111101;
    krom[773] = 9'b110111100;
    krom[774] = 9'b100111100;
    krom[775] = 9'b111111100;
    krom[777] = 9'b111011100;
    krom[778] = 9'b101011100;
    krom[779] = 9'b100011100;
    krom[780] = 9'b101111100;
    krom[781] = 9'b110011100;
    krom[786] = 9'b110000011;
    krom[787] = 9'b101100011;
    krom[788] = 9'b100000011;
    krom[789] = 9'b101000011;
    krom[790] = 9'b111000011;
    krom[791] = 9'b011100011;
    krom[792] = 9'b111100011;
    krom[793] = 9'b100100011;
    krom[794] = 9'b110100011;
    krom[795] = 9'b000000011;
    krom[796] = 9'b001100011;
    krom[797] = 9'b010000011;
    krom[802] = 9'b110010011;
    krom[803] = 9'b101110011;
    krom[804] = 9'b100010011;
    krom[805] = 9'b101010011;
    krom[806] = 9'b111010011;
    krom[807] = 9'b011110011;
    krom[808] = 9'b111110011;
    krom[809] = 9'b100110011;
    krom[810] = 9'b110110011;
    krom[811] = 9'b000010011;
    krom[812] = 9'b001110011;
    krom[813] = 9'b010010011;
    krom[818] = 9'b010011000;
    krom[819] = 9'b001111000;
    krom[820] = 9'b000011000;
    krom[821] = 9'b001011000;
    krom[822] = 9'b011011000;
    krom[824] = 9'b011111000;
    krom[825] = 9'b000111000;
    krom[826] = 9'b010111000;
    krom[834] = 9'b110001011;
    krom[835] = 9'b101101011;
    krom[836] = 9'b100001011;
    krom[837] = 9'b101001011;
    krom[838] = 9'b111001011;
    krom[839] = 9'b011101011;
    krom[840] = 9'b111101011;
    krom[841] = 9'b100101011;
    krom[842] = 9'b110101011;
    krom[843] = 9'b000001011;
    krom[844] = 9'b001101011;
    krom[845] = 9'b010001011;
    krom[850] = 9'b010000100;
    krom[851] = 9'b001100100;
    krom[852] = 9'b000000100;
    krom[853] = 9'b001000100;
    krom[854] = 9'b011000100;
    krom[856] = 9'b011100100;
    krom[857] = 9'b000100100;
    krom[858] = 9'b010100100;
    krom[866] = 9'b010011011;
    krom[867] = 9'b001111011;
    krom[868] = 9'b000011011;
    krom[869] = 9'b001011011;
    krom[870] = 9'b011011011;
    krom[872] = 9'b011111011;
    krom[873] = 9'b000111011;
    krom[874] = 9'b010111011;
    krom[901] = 9'b010100111;
    krom[902] = 9'b000100111;
    krom[903] = 9'b011100111;
    krom[905] = 9'b011000111;
    krom[906] = 9'b001000111;
    krom[907] = 9'b000000111;
    krom[908] = 9'b001100111;
    krom[909] = 9'b010000111;
    krom[914] = 9'b010001000;
    krom[915] = 9'b001101000;
    krom[916] = 9'b000001000;
    krom[917] = 9'b001001000;
    krom[918] = 9'b011001000;
    krom[920] = 9'b011101000;
    krom[921] = 9'b000101000;
    krom[922] = 9'b010101000;
    krom[930] = 9'b010010111;
    krom[931] = 9'b001110111;
    krom[932] = 9'b000010111;
    krom[933] = 9'b001010111;
    krom[934] = 9'b011010111;
    krom[936] = 9'b011110111;
    krom[937] = 9'b000110111;
    krom[938] = 9'b010110111;
  end

  initial begin
    drom[85] = 9'b101010111;
    drom[86] = 9'b111010111;
    drom[89] = 9'b100110111;
    drom[90] = 9'b110110111;
    drom[91] = 9'b100010111;
    drom[92] = 9'b101110111;
    drom[93] = 9'b110010111;
    drom[94] = 9'b111110111;
    drom[101] = 9'b101001000;
    drom[102] = 9'b111001000;
    drom[105] = 9'b100101000;
    drom[106] = 9'b110101000;
    drom[107] = 9'b100001000;
    drom[108] = 9'b101101000;
    drom[109] = 9'b110001000;
    drom[110] = 9'b111101000;
    drom[113] = 9'b111100111;
    drom[114] = 9'b110000111;
    drom[115] = 9'b101100111;
    drom[116] = 9'b100000111;
    drom[117] = 9'b101000111;
    drom[118] = 9'b111000111;
    drom[121] = 9'b100100111;
    drom[122] = 9'b110100111;
    drom[149] = 9'b101011011;
    drom[150] = 9'b111011011;
    drom[153] = 9'b100111011;
    drom[154] = 9'b110111011;
    drom[155] = 9'b100011011;
    drom[156] = 9'b101111011;
    drom[157] = 9'b110011011;
    drom[158] = 9'b111111011;
    drom[165] = 9'b101000100;
    drom[166] = 9'b111000100;
    drom[169] = 9'b100100100;
    drom[170] = 9'b110100100;
    drom[171] = 9'b100000100;
    drom[172] = 9'b101100100;
    drom[173] = 9'b110000100;
    drom[174] = 9'b111100100;
    drom[177] = 9'b111110100;
    drom[178] = 9'b110010100;
    drom[179] = 9'b101110100;
    drom[180] = 9'b100010100;
    drom[181] = 9'b101010100;
    drom[182] = 9'b111010100;
    drom[183] = 9'b011110100;
    drom[185] = 9'b100110100;
    drom[186] = 9'b110110100;
    drom[187] = 9'b000010100;
    drom[188] = 9'b001110100;
    drom[189] = 9'b010010100;
    drom[197] = 9'b101011000;
    drom[198] = 9'b111011000;
    drom[201] = 9'b100111000;
    drom[202] = 9'b110111000;
    drom[203] = 9'b100011000;
    drom[204] = 9'b101111000;
    drom[205] = 9'b110011000;
    drom[206] = 9'b111111000;
    drom[209] = 9'b111101100;
    drom[210] = 9'b110001100;
    drom[211] = 9'b101101100;
    drom[212] = 9'b100001100;
    drom[213] = 9'b101001100;
    drom[214] = 9'b111001100;
    drom[217] = 9'b100101100;
    drom[218] = 9'b110101100;
    drom[219] = 9'b000001100;
    drom[220] = 9'b001101100;
    drom[221] = 9'b010001100;
    drom[222] = 9'b011101100;
    drom[225] = 9'b111111100;
    drom[226] = 9'b110011100;
    drom[227] = 9'b101111100;
    drom[228] = 9'b100011100;
    drom[229] = 9'b101011100;
    drom[230] = 9'b111011100;
    drom[233] = 9'b100111100;
    drom[234] = 9'b110111100;
    drom[235] = 9'b000011100;
    drom[236] = 9'b001111100;
    drom[237] = 9'b010011100;
    drom[238] = 9'b011111100;
    drom[277] = 9'b101011101;
    drom[278] = 9'b111011101;
    drom[281] = 9'b100111101;
    drom[282] = 9'b110111101;
    drom[283] = 9'b100011101;
    drom[284] = 9'b101111101;
    drom[285] = 9'b110011101;
    drom[286] = 9'b111111101;
    drom[293] = 9'b101000010;
    drom[294] = 9'b111000010;
    drom[297] = 9'b100100010;
    drom[298] = 9'b110100010;
    drom[299] = 9'b100000010;
    drom[300] = 9'b101100010;
    drom[301] = 9'b110000010;
    drom[302] = 9'b111100010;
    drom[305] = 9'b111110010;
    drom[306] = 9'b110010010;
    drom[307] = 9'b101110010;
    drom[308] = 9'b100010010;
    drom[309] = 9'b101010010;
    drom[310] = 9'b111010010;
    drom[311] = 9'b011110010;
    drom[313] = 9'b100110010;
    drom[314] = 9'b110110010;
    drom[315] = 9'b000010010;
    drom[316] = 9'b001110010;
    drom[317] = 9'b010010010;
    drom[325] = 9'b101011111;
    drom[326] = 9'b111011111;
    drom[329] = 9'b100111111;
    drom[330] = 9'b110111111;
    drom[331] = 9'b100011111;
    drom[332] = 9'b101111111;
    drom[333] = 9'b110011111;
    drom[334] = 9'b111111111;
    drom[337] = 9'b111101010;
    drom[338] = 9'b110001010;
    drom[339] = 9'b101101010;
    drom[340] = 9'b100001010;
    drom[341] = 9'b101001010;
    drom[342] = 9'b111001010;
    drom[345] = 9'b100101010;
    drom[346] = 9'b110101010;
    drom[347] = 9'b000001010;
    drom[348] = 9'b001101010;
    drom[349] = 9'b010001010;
    drom[350] = 9'b011101010;
    drom[353] = 9'b111111010;
    drom[354] = 9'b110011010;
    drom[355] = 9'b101111010;
    drom[356] = 9'b100011010;
    drom[357] = 9'b101011010;
    drom[358] = 9'b111011010;
    drom[361] = 9'b100111010;
    drom[362] = 9'b110111010;
    drom[363] = 9'b000011010;
    drom[364] = 9'b001111010;
    drom[365] = 9'b010011010;
    drom[366] = 9'b011111010;
    drom[369] = 9'b011101111;
    drom[370] = 9'b010001111;
    drom[371] = 9'b001101111;
    drom[372] = 9'b000001111;
    drom[373] = 9'b001001111;
    drom[374] = 9'b011001111;
    drom[377] = 9'b000101111;
    drom[378] = 9'b010101111;
    drom[389] = 9'b101000000;
    drom[390] = 9'b111000000;
    drom[393] = 9'b100100000;
    drom[394] = 9'b110100000;
    drom[395] = 9'b100000000;
    drom[396] = 9'b101100000;
    drom[397] = 9'b110000000;
    drom[398] = 9'b111100000;
    drom[401] = 9'b111100110;
    drom[402] = 9'b110000110;
    drom[403] = 9'b101100110;
    drom[404] = 9'b100000110;
    drom[405] = 9'b101000110;
    drom[406] = 9'b111000110;
    drom[409] = 9'b100100110;
    drom[410] = 9'b110100110;
    drom[411] = 9'b000000110;
    drom[412] = 9'b001100110;
    drom[413] = 9'b010000110;
    drom[414] = 9'b011100110;
    drom[417] = 9'b111110110;
    drom[418] = 9'b110010110;
    drom[419] = 9'b101110110;
    drom[420] = 9'b100010110;
    drom[421] = 9'b101010110;
    drom[422] = 9'b111010110;
    drom[425] = 9'b100110110;
    drom[426] = 9'b110110110;
    drom[427] = 9'b000010110;
    drom[428] = 9'b001110110;
    drom[429] = 9'b010010110;
    drom[430] = 9'b011110110;
    drom[433] = 9'b011110000;
    drom[434] = 9'b010010000;
    drom[435] = 9'b001110000;
    drom[436] = 9'b000010000;
    drom[437] = 9'b001010000;
    drom[438] = 9'b011010000;
    drom[441] = 9'b000110000;
    drom[442] = 9'b010110000;
    drom[450] = 9'b110001110;
    drom[451] = 9'b101101110;
    drom[452] = 9'b100001110;
    drom[453] = 9'b101001110;
    drom[454] = 9'b111001110;
    drom[456] = 9'b111101110;
    drom[457] = 9'b100101110;
    drom[458] = 9'b110101110;
    drom[459] = 9'b000001110;
    drom[460] = 9'b001101110;
    drom[461] = 9'b010001110;
    drom[462] = 9'b011101110;
    drom[465] = 9'b011100001;
    drom[466] = 9'b010000001;
    drom[467] = 9'b001100001;
    drom[468] = 9'b000000001;
    drom[469] = 9'b001000001;
    drom[470] = 9'b011000001;
    drom[473] = 9'b000100001;
    drom[474] = 9'b010100001;
    drom[481] = 9'b011111110;
    drom[482] = 9'b010011110;
    drom[483] = 9'b001111110;
    drom[484] = 9'b000011110;
    drom[485] = 9'b001011110;
    drom[486] = 9'b011011110;
    drom[489] = 9'b000111110;
    drom[490] = 9'b010111110;
    drom[533] = 9'b101011110;
    drom[534] = 9'b111011110;
    drom[537] = 9'b100111110;
    drom[538] = 9'b110111110;
    drom[539] = 9'b100011110;
    drom[540] = 9'b101111110;
    drom[541] = 9'b110011110;
    drom[542] = 9'b111111110;
    drom[549] = 9'b101000001;
    drom[550] = 9'b111000001;
    drom[553] = 9'b100100001;
    drom[554] = 9'b110100001;
    drom[555] = 9'b100000001;
    drom[556] = 9'b101100001;
    drom[557] = 9'b110000001;
    drom[558] = 9'b111100001;
    drom[561] = 9'b111110001;
    drom[562] = 9'b110010001;
    drom[563] = 9'b101110001;
    drom[564] = 9'b100010001;
    drom[565] = 9'b101010001;
    drom[566] = 9'b111010001;
    drom[567] = 9'b011110001;
    drom[569] = 9'b100110001;
    drom[570] = 9'b110110001;
    drom[571] = 9'b000010001;
    drom[572] = 9'b001110001;
    drom[573] = 9'b010010001;
    drom[581] = 9'b101010000;
    drom[582] = 9'b111010000;
    drom[585] = 9'b100110000;
    drom[586] = 9'b110110000;
    drom[587] = 9'b100010000;
    drom[588] = 9'b101110000;
    drom[589] = 9'b110010000;
    drom[590] = 9'b111110000;
    drom[593] = 9'b111101001;
    drom[594] = 9'b110001001;
    drom[595] = 9'b101101001;
    drom[596] = 9'b100001001;
    drom[597] = 9'b101001001;
    drom[598] = 9'b111001001;
    drom[601] = 9'b100101001;
    drom[602] = 9'b110101001;
    drom[603] = 9'b000001001;
    drom[604] = 9'b001101001;
    drom[605] = 9'b010001001;
    drom[606] = 9'b011101001;
    drom[609] = 9'b111111001;
    drom[610] = 9'b110011001;
    drom[611] = 9'b101111001;
    drom[612] = 9'b100011001;
    drom[613] = 9'b101011001;
    drom[614] = 9'b111011001;
    drom[617] = 9'b100111001;
    drom[618] = 9'b110111001;
    drom[619] = 9'b000011001;
    drom[620] = 9'b001111001;
    drom[621] = 9'b010011001;
    drom[622] = 9'b011111001;
    drom[625] = 9'b011100000;
    drom[626] = 9'b010000000;
    drom[627] = 9'b001100000;
    drom[628] = 9'b000000000;
    drom[629] = 9'b001000000;
    drom[630] = 9'b011000000;
    drom[633] = 9'b000100000;
    drom[634] = 9'b010100000;
    drom[645] = 9'b101001111;
    drom[646] = 9'b111001111;
    drom[649] = 9'b100101111;
    drom[650] = 9'b110101111;
    drom[651] = 9'b100001111;
    drom[652] = 9'b101101111;
    drom[653] = 9'b110001111;
    drom[654] = 9'b111101111;
    drom[657] = 9'b111100101;
    drom[658] = 9'b110000101;
    drom[659] = 9'b101100101;
    drom[660] = 9'b100000101;
    drom[661] = 9'b101000101;
    drom[662] = 9'b111000101;
    drom[665] = 9'b100100101;
    drom[666] = 9'b110100101;
    drom[667] = 9'b000000101;
    drom[668] = 9'b001100101;
    drom[669] = 9'b010000101;
    drom[670] = 9'b011100101;
    drom[673] = 9'b111110101;
    drom[674] = 9'b110010101;
    drom[675] = 9'b101110101;
    drom[676] = 9'b100010101;
    drom[677] = 9'b101010101;
    drom[678] = 9'b111010101;
    drom[681] = 9'b100110101;
    drom[682] = 9'b110110101;
    drom[683] = 9'b000010101;
    drom[684] = 9'b001110101;
    drom[685] = 9'b010010101;
    drom[686] = 9'b011110101;
    drom[689] = 9'b011111111;
    drom[690] = 9'b010011111;
    drom[691] = 9'b001111111;
    drom[692] = 9'b000011111;
    drom[693] = 9'b001011111;
    drom[694] = 9'b011011111;
    drom[697] = 9'b000111111;
    drom[698] = 9'b010111111;
    drom[706] = 9'b110001101;
    drom[707] = 9'b101101101;
    drom[708] = 9'b100001101;
    drom[709] = 9'b101001101;
    drom[710] = 9'b111001101;
    drom[712] = 9'b111101101;
    drom[713] = 9'b100101101;
    drom[714] = 9'b110101101;
    drom[715] = 9'b000001101;
    drom[716] = 9'b001101101;
    drom[717] = 9'b010001101;
    drom[718] = 9'b011101101;
    drom[721] = 9'b011100010;
    drom[722] = 9'b010000010;
    drom[723] = 9'b001100010;
    drom[724] = 9'b000000010;
    drom[725] = 9'b001000010;
    drom[726] = 9'b011000010;
    drom[729] = 9'b000100010;
    drom[730] = 9'b010100010;
    drom[737] = 9'b011111101;
    drom[738] = 9'b010011101;
    drom[739] = 9'b001111101;
    drom[740] = 9'b000011101;
    drom[741] = 9'b001011101;
    drom[742] = 9'b011011101;
    drom[745] = 9'b000111101;
    drom[746] = 9'b010111101;
    drom[785] = 9'b111100011;
    drom[786] = 9'b110000011;
    drom[787] = 9'b101100011;
    drom[788] = 9'b100000011;
    drom[789] = 9'b101000011;
    drom[790] = 9'b111000011;
    drom[793] = 9'b100100011;
    drom[794] = 9'b110100011;
    drom[795] = 9'b000000011;
    drom[796] = 9'b001100011;
    drom[797] = 9'b010000011;
    drom[798] = 9'b011100011;
    drom[801] = 9'b111110011;
    drom[802] = 9'b110010011;
    drom[803] = 9'b101110011;
    drom[804] = 9'b100010011;
    drom[805] = 9'b101010011;
    drom[806] = 9'b111010011;
    drom[809] = 9'b100110011;
    drom[810] = 9'b110110011;
    drom[811] = 9'b000010011;
    drom[812] = 9'b001110011;
    drom[813] = 9'b010010011;
    drom[814] = 9'b011110011;
    drom[817] = 9'b011111000;
    drom[818] = 9'b010011000;
    drom[819] = 9'b001111000;
    drom[820] = 9'b000011000;
    drom[821] = 9'b001011000;
    drom[822] = 9'b011011000;
    drom[825] = 9'b000111000;
    drom[826] = 9'b010111000;
    drom[834] = 9'b110001011;
    drom[835] = 9'b101101011;
    drom[836] = 9'b100001011;
    drom[837] = 9'b101001011;
    drom[838] = 9'b111001011;
    drom[840] = 9'b111101011;
    drom[841] = 9'b100101011;
    drom[842] = 9'b110101011;
    drom[843] = 9'b000001011;
    drom[844] = 9'b001101011;
    drom[845] = 9'b010001011;
    drom[846] = 9'b011101011;
    drom[849] = 9'b011100100;
    drom[850] = 9'b010000100;
    drom[851] = 9'b001100100;
    drom[852] = 9'b000000100;
    drom[853] = 9'b001000100;
    drom[854] = 9'b011000100;
    drom[857] = 9'b000100100;
    drom[858] = 9'b010100100;
    drom[865] = 9'b011111011;
    drom[866] = 9'b010011011;
    drom[867] = 9'b001111011;
    drom[868] = 9'b000011011;
    drom[869] = 9'b001011011;
    drom[870] = 9'b011011011;
    drom[873] = 9'b000111011;
    drom[874] = 9'b010111011;
    drom[901] = 9'b001000111;
    drom[902] = 9'b011000111;
    drom[905] = 9'b000100111;
    drom[906] = 9'b010100111;
    drom[907] = 9'b000000111;
    drom[908] = 9'b001100111;
    drom[909] = 9'b010000111;
    drom[910] = 9'b011100111;
    drom[913] = 9'b011101000;
    drom[914] = 9'b010001000;
    drom[915] = 9'b001101000;
    drom[916] = 9'b000001000;
    drom[917] = 9'b001001000;
    drom[918] = 9'b011001000;
    drom[921] = 9'b000101000;
    drom[922] = 9'b010101000;
    drom[929] = 9'b011110111;
    drom[930] = 9'b010010111;
    drom[931] = 9'b001110111;
    drom[932] = 9'b000010111;
    drom[933] = 9'b001010111;
    drom[934] = 9'b011010111;
    drom[937] = 9'b000110111;
    drom[938] = 9'b010110111;
  end

endmodule : decoder_8b10b
