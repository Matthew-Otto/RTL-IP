// encodes bytes and control symbols to 8b/10b scheme
// outputs data in the order abcdei fghj
// 10b symbols should be serialized MSB first

module encoder_8b10b (
  input  logic       clk,
  input  logic       reset,
  input  logic       input_valid,
  input  logic       input_ctrl,
  input  logic [7:0] input_data,
  output logic [9:0] output_data
);

  logic        rd, next_rd;
  logic [9:0]  rom_addr;
  logic [10:0] rom_read;

  always_ff @(posedge clk)
    if (reset)            rd <= 0;
    else if (input_valid) rd <= next_rd;

  assign rom_addr = {input_ctrl,rd,input_data};
  assign rom_read = rom[rom_addr];
  assign output_data = rom_read[9:0];
  assign next_rd = rom_read[10];
  
  logic [10:0] rom [1023:0];
  
  initial begin
    rom[0] = 11'b01001110100;	// -D00.0-
    rom[1] = 11'b00111010100;	// -D01.0-
    rom[2] = 11'b01011010100;	// -D02.0-
    rom[3] = 11'b11100011011;	// -D03.0+
    rom[4] = 11'b01101010100;	// -D04.0-
    rom[5] = 11'b11010011011;	// -D05.0+
    rom[6] = 11'b10110011011;	// -D06.0+
    rom[7] = 11'b11110001011;	// -D07.0+
    rom[8] = 11'b01110010100;	// -D08.0-
    rom[9] = 11'b11001011011;	// -D09.0+
    rom[10] = 11'b10101011011;	// -D10.0+
    rom[11] = 11'b11101001011;	// -D11.0+
    rom[12] = 11'b10011011011;	// -D12.0+
    rom[13] = 11'b11011001011;	// -D13.0+
    rom[14] = 11'b10111001011;	// -D14.0+
    rom[15] = 11'b00101110100;	// -D15.0-
    rom[16] = 11'b00110110100;	// -D16.0-
    rom[17] = 11'b11000111011;	// -D17.0+
    rom[18] = 11'b10100111011;	// -D18.0+
    rom[19] = 11'b11100101011;	// -D19.0+
    rom[20] = 11'b10010111011;	// -D20.0+
    rom[21] = 11'b11010101011;	// -D21.0+
    rom[22] = 11'b10110101011;	// -D22.0+
    rom[23] = 11'b01110100100;	// -D23.0-
    rom[24] = 11'b01100110100;	// -D24.0-
    rom[25] = 11'b11001101011;	// -D25.0+
    rom[26] = 11'b10101101011;	// -D26.0+
    rom[27] = 11'b01101100100;	// -D27.0-
    rom[28] = 11'b10011101011;	// -D28.0+
    rom[29] = 11'b01011100100;	// -D29.0-
    rom[30] = 11'b00111100100;	// -D30.0-
    rom[31] = 11'b01010110100;	// -D31.0-
    rom[32] = 11'b11001111001;	// -D00.1+
    rom[33] = 11'b10111011001;	// -D01.1+
    rom[34] = 11'b11011011001;	// -D02.1+
    rom[35] = 11'b01100011001;	// -D03.1-
    rom[36] = 11'b11101011001;	// -D04.1+
    rom[37] = 11'b01010011001;	// -D05.1-
    rom[38] = 11'b00110011001;	// -D06.1-
    rom[39] = 11'b01110001001;	// -D07.1-
    rom[40] = 11'b11110011001;	// -D08.1+
    rom[41] = 11'b01001011001;	// -D09.1-
    rom[42] = 11'b00101011001;	// -D10.1-
    rom[43] = 11'b01101001001;	// -D11.1-
    rom[44] = 11'b00011011001;	// -D12.1-
    rom[45] = 11'b01011001001;	// -D13.1-
    rom[46] = 11'b00111001001;	// -D14.1-
    rom[47] = 11'b10101111001;	// -D15.1+
    rom[48] = 11'b10110111001;	// -D16.1+
    rom[49] = 11'b01000111001;	// -D17.1-
    rom[50] = 11'b00100111001;	// -D18.1-
    rom[51] = 11'b01100101001;	// -D19.1-
    rom[52] = 11'b00010111001;	// -D20.1-
    rom[53] = 11'b01010101001;	// -D21.1-
    rom[54] = 11'b00110101001;	// -D22.1-
    rom[55] = 11'b11110101001;	// -D23.1+
    rom[56] = 11'b11100111001;	// -D24.1+
    rom[57] = 11'b01001101001;	// -D25.1-
    rom[58] = 11'b00101101001;	// -D26.1-
    rom[59] = 11'b11101101001;	// -D27.1+
    rom[60] = 11'b00011101001;	// -D28.1-
    rom[61] = 11'b11011101001;	// -D29.1+
    rom[62] = 11'b10111101001;	// -D30.1+
    rom[63] = 11'b11010111001;	// -D31.1+
    rom[64] = 11'b11001110101;	// -D00.2+
    rom[65] = 11'b10111010101;	// -D01.2+
    rom[66] = 11'b11011010101;	// -D02.2+
    rom[67] = 11'b01100010101;	// -D03.2-
    rom[68] = 11'b11101010101;	// -D04.2+
    rom[69] = 11'b01010010101;	// -D05.2-
    rom[70] = 11'b00110010101;	// -D06.2-
    rom[71] = 11'b01110000101;	// -D07.2-
    rom[72] = 11'b11110010101;	// -D08.2+
    rom[73] = 11'b01001010101;	// -D09.2-
    rom[74] = 11'b00101010101;	// -D10.2-
    rom[75] = 11'b01101000101;	// -D11.2-
    rom[76] = 11'b00011010101;	// -D12.2-
    rom[77] = 11'b01011000101;	// -D13.2-
    rom[78] = 11'b00111000101;	// -D14.2-
    rom[79] = 11'b10101110101;	// -D15.2+
    rom[80] = 11'b10110110101;	// -D16.2+
    rom[81] = 11'b01000110101;	// -D17.2-
    rom[82] = 11'b00100110101;	// -D18.2-
    rom[83] = 11'b01100100101;	// -D19.2-
    rom[84] = 11'b00010110101;	// -D20.2-
    rom[85] = 11'b01010100101;	// -D21.2-
    rom[86] = 11'b00110100101;	// -D22.2-
    rom[87] = 11'b11110100101;	// -D23.2+
    rom[88] = 11'b11100110101;	// -D24.2+
    rom[89] = 11'b01001100101;	// -D25.2-
    rom[90] = 11'b00101100101;	// -D26.2-
    rom[91] = 11'b11101100101;	// -D27.2+
    rom[92] = 11'b00011100101;	// -D28.2-
    rom[93] = 11'b11011100101;	// -D29.2+
    rom[94] = 11'b10111100101;	// -D30.2+
    rom[95] = 11'b11010110101;	// -D31.2+
    rom[96] = 11'b11001110011;	// -D00.3+
    rom[97] = 11'b10111010011;	// -D01.3+
    rom[98] = 11'b11011010011;	// -D02.3+
    rom[99] = 11'b01100011100;	// -D03.3-
    rom[100] = 11'b11101010011;	// -D04.3+
    rom[101] = 11'b01010011100;	// -D05.3-
    rom[102] = 11'b00110011100;	// -D06.3-
    rom[103] = 11'b01110001100;	// -D07.3-
    rom[104] = 11'b11110010011;	// -D08.3+
    rom[105] = 11'b01001011100;	// -D09.3-
    rom[106] = 11'b00101011100;	// -D10.3-
    rom[107] = 11'b01101001100;	// -D11.3-
    rom[108] = 11'b00011011100;	// -D12.3-
    rom[109] = 11'b01011001100;	// -D13.3-
    rom[110] = 11'b00111001100;	// -D14.3-
    rom[111] = 11'b10101110011;	// -D15.3+
    rom[112] = 11'b10110110011;	// -D16.3+
    rom[113] = 11'b01000111100;	// -D17.3-
    rom[114] = 11'b00100111100;	// -D18.3-
    rom[115] = 11'b01100101100;	// -D19.3-
    rom[116] = 11'b00010111100;	// -D20.3-
    rom[117] = 11'b01010101100;	// -D21.3-
    rom[118] = 11'b00110101100;	// -D22.3-
    rom[119] = 11'b11110100011;	// -D23.3+
    rom[120] = 11'b11100110011;	// -D24.3+
    rom[121] = 11'b01001101100;	// -D25.3-
    rom[122] = 11'b00101101100;	// -D26.3-
    rom[123] = 11'b11101100011;	// -D27.3+
    rom[124] = 11'b00011101100;	// -D28.3-
    rom[125] = 11'b11011100011;	// -D29.3+
    rom[126] = 11'b10111100011;	// -D30.3+
    rom[127] = 11'b11010110011;	// -D31.3+
    rom[128] = 11'b01001110010;	// -D00.4-
    rom[129] = 11'b00111010010;	// -D01.4-
    rom[130] = 11'b01011010010;	// -D02.4-
    rom[131] = 11'b11100011101;	// -D03.4+
    rom[132] = 11'b01101010010;	// -D04.4-
    rom[133] = 11'b11010011101;	// -D05.4+
    rom[134] = 11'b10110011101;	// -D06.4+
    rom[135] = 11'b11110001101;	// -D07.4+
    rom[136] = 11'b01110010010;	// -D08.4-
    rom[137] = 11'b11001011101;	// -D09.4+
    rom[138] = 11'b10101011101;	// -D10.4+
    rom[139] = 11'b11101001101;	// -D11.4+
    rom[140] = 11'b10011011101;	// -D12.4+
    rom[141] = 11'b11011001101;	// -D13.4+
    rom[142] = 11'b10111001101;	// -D14.4+
    rom[143] = 11'b00101110010;	// -D15.4-
    rom[144] = 11'b00110110010;	// -D16.4-
    rom[145] = 11'b11000111101;	// -D17.4+
    rom[146] = 11'b10100111101;	// -D18.4+
    rom[147] = 11'b11100101101;	// -D19.4+
    rom[148] = 11'b10010111101;	// -D20.4+
    rom[149] = 11'b11010101101;	// -D21.4+
    rom[150] = 11'b10110101101;	// -D22.4+
    rom[151] = 11'b01110100010;	// -D23.4-
    rom[152] = 11'b01100110010;	// -D24.4-
    rom[153] = 11'b11001101101;	// -D25.4+
    rom[154] = 11'b10101101101;	// -D26.4+
    rom[155] = 11'b01101100010;	// -D27.4-
    rom[156] = 11'b10011101101;	// -D28.4+
    rom[157] = 11'b01011100010;	// -D29.4-
    rom[158] = 11'b00111100010;	// -D30.4-
    rom[159] = 11'b01010110010;	// -D31.4-
    rom[160] = 11'b11001111010;	// -D00.5+
    rom[161] = 11'b10111011010;	// -D01.5+
    rom[162] = 11'b11011011010;	// -D02.5+
    rom[163] = 11'b01100011010;	// -D03.5-
    rom[164] = 11'b11101011010;	// -D04.5+
    rom[165] = 11'b01010011010;	// -D05.5-
    rom[166] = 11'b00110011010;	// -D06.5-
    rom[167] = 11'b01110001010;	// -D07.5-
    rom[168] = 11'b11110011010;	// -D08.5+
    rom[169] = 11'b01001011010;	// -D09.5-
    rom[170] = 11'b00101011010;	// -D10.5-
    rom[171] = 11'b01101001010;	// -D11.5-
    rom[172] = 11'b00011011010;	// -D12.5-
    rom[173] = 11'b01011001010;	// -D13.5-
    rom[174] = 11'b00111001010;	// -D14.5-
    rom[175] = 11'b10101111010;	// -D15.5+
    rom[176] = 11'b10110111010;	// -D16.5+
    rom[177] = 11'b01000111010;	// -D17.5-
    rom[178] = 11'b00100111010;	// -D18.5-
    rom[179] = 11'b01100101010;	// -D19.5-
    rom[180] = 11'b00010111010;	// -D20.5-
    rom[181] = 11'b01010101010;	// -D21.5-
    rom[182] = 11'b00110101010;	// -D22.5-
    rom[183] = 11'b11110101010;	// -D23.5+
    rom[184] = 11'b11100111010;	// -D24.5+
    rom[185] = 11'b01001101010;	// -D25.5-
    rom[186] = 11'b00101101010;	// -D26.5-
    rom[187] = 11'b11101101010;	// -D27.5+
    rom[188] = 11'b00011101010;	// -D28.5-
    rom[189] = 11'b11011101010;	// -D29.5+
    rom[190] = 11'b10111101010;	// -D30.5+
    rom[191] = 11'b11010111010;	// -D31.5+
    rom[192] = 11'b11001110110;	// -D00.6+
    rom[193] = 11'b10111010110;	// -D01.6+
    rom[194] = 11'b11011010110;	// -D02.6+
    rom[195] = 11'b01100010110;	// -D03.6-
    rom[196] = 11'b11101010110;	// -D04.6+
    rom[197] = 11'b01010010110;	// -D05.6-
    rom[198] = 11'b00110010110;	// -D06.6-
    rom[199] = 11'b01110000110;	// -D07.6-
    rom[200] = 11'b11110010110;	// -D08.6+
    rom[201] = 11'b01001010110;	// -D09.6-
    rom[202] = 11'b00101010110;	// -D10.6-
    rom[203] = 11'b01101000110;	// -D11.6-
    rom[204] = 11'b00011010110;	// -D12.6-
    rom[205] = 11'b01011000110;	// -D13.6-
    rom[206] = 11'b00111000110;	// -D14.6-
    rom[207] = 11'b10101110110;	// -D15.6+
    rom[208] = 11'b10110110110;	// -D16.6+
    rom[209] = 11'b01000110110;	// -D17.6-
    rom[210] = 11'b00100110110;	// -D18.6-
    rom[211] = 11'b01100100110;	// -D19.6-
    rom[212] = 11'b00010110110;	// -D20.6-
    rom[213] = 11'b01010100110;	// -D21.6-
    rom[214] = 11'b00110100110;	// -D22.6-
    rom[215] = 11'b11110100110;	// -D23.6+
    rom[216] = 11'b11100110110;	// -D24.6+
    rom[217] = 11'b01001100110;	// -D25.6-
    rom[218] = 11'b00101100110;	// -D26.6-
    rom[219] = 11'b11101100110;	// -D27.6+
    rom[220] = 11'b00011100110;	// -D28.6-
    rom[221] = 11'b11011100110;	// -D29.6+
    rom[222] = 11'b10111100110;	// -D30.6+
    rom[223] = 11'b11010110110;	// -D31.6+
    rom[224] = 11'b01001110001;	// -D00.7-
    rom[225] = 11'b00111010001;	// -D01.7-
    rom[226] = 11'b01011010001;	// -D02.7-
    rom[227] = 11'b11100011110;	// -D03.7+
    rom[228] = 11'b01101010001;	// -D04.7-
    rom[229] = 11'b11010011110;	// -D05.7+
    rom[230] = 11'b10110011110;	// -D06.7+
    rom[231] = 11'b11110001110;	// -D07.7+
    rom[232] = 11'b01110010001;	// -D08.7-
    rom[233] = 11'b11001011110;	// -D09.7+
    rom[234] = 11'b10101011110;	// -D10.7+
    rom[235] = 11'b11101001110;	// -D11.7+
    rom[236] = 11'b10011011110;	// -D12.7+
    rom[237] = 11'b11011001110;	// -D13.7+
    rom[238] = 11'b10111001110;	// -D14.7+
    rom[239] = 11'b00101110001;	// -D15.7-
    rom[240] = 11'b00110110001;	// -D16.7-
    rom[241] = 11'b11000110111;	// -D17.7+
    rom[242] = 11'b10100110111;	// -D18.7+
    rom[243] = 11'b11100101110;	// -D19.7+
    rom[244] = 11'b10010110111;	// -D20.7+
    rom[245] = 11'b11010101110;	// -D21.7+
    rom[246] = 11'b10110101110;	// -D22.7+
    rom[247] = 11'b01110100001;	// -D23.7-
    rom[248] = 11'b01100110001;	// -D24.7-
    rom[249] = 11'b11001101110;	// -D25.7+
    rom[250] = 11'b10101101110;	// -D26.7+
    rom[251] = 11'b01101100001;	// -D27.7-
    rom[252] = 11'b10011101110;	// -D28.7+
    rom[253] = 11'b01011100001;	// -D29.7-
    rom[254] = 11'b00111100001;	// -D30.7-
    rom[255] = 11'b01010110001;	// -D31.7-
    rom[256] = 11'b10110001011;	// +D00.0+
    rom[257] = 11'b11000101011;	// +D01.0+
    rom[258] = 11'b10100101011;	// +D02.0+
    rom[259] = 11'b01100010100;	// +D03.0-
    rom[260] = 11'b10010101011;	// +D04.0+
    rom[261] = 11'b01010010100;	// +D05.0-
    rom[262] = 11'b00110010100;	// +D06.0-
    rom[263] = 11'b00001110100;	// +D07.0-
    rom[264] = 11'b10001101011;	// +D08.0+
    rom[265] = 11'b01001010100;	// +D09.0-
    rom[266] = 11'b00101010100;	// +D10.0-
    rom[267] = 11'b01101000100;	// +D11.0-
    rom[268] = 11'b00011010100;	// +D12.0-
    rom[269] = 11'b01011000100;	// +D13.0-
    rom[270] = 11'b00111000100;	// +D14.0-
    rom[271] = 11'b11010001011;	// +D15.0+
    rom[272] = 11'b11001001011;	// +D16.0+
    rom[273] = 11'b01000110100;	// +D17.0-
    rom[274] = 11'b00100110100;	// +D18.0-
    rom[275] = 11'b01100100100;	// +D19.0-
    rom[276] = 11'b00010110100;	// +D20.0-
    rom[277] = 11'b01010100100;	// +D21.0-
    rom[278] = 11'b00110100100;	// +D22.0-
    rom[279] = 11'b10001011011;	// +D23.0+
    rom[280] = 11'b10011001011;	// +D24.0+
    rom[281] = 11'b01001100100;	// +D25.0-
    rom[282] = 11'b00101100100;	// +D26.0-
    rom[283] = 11'b10010011011;	// +D27.0+
    rom[284] = 11'b00011100100;	// +D28.0-
    rom[285] = 11'b10100011011;	// +D29.0+
    rom[286] = 11'b11000011011;	// +D30.0+
    rom[287] = 11'b10101001011;	// +D31.0+
    rom[288] = 11'b00110001001;	// +D00.1-
    rom[289] = 11'b01000101001;	// +D01.1-
    rom[290] = 11'b00100101001;	// +D02.1-
    rom[291] = 11'b11100011001;	// +D03.1+
    rom[292] = 11'b00010101001;	// +D04.1-
    rom[293] = 11'b11010011001;	// +D05.1+
    rom[294] = 11'b10110011001;	// +D06.1+
    rom[295] = 11'b10001111001;	// +D07.1+
    rom[296] = 11'b00001101001;	// +D08.1-
    rom[297] = 11'b11001011001;	// +D09.1+
    rom[298] = 11'b10101011001;	// +D10.1+
    rom[299] = 11'b11101001001;	// +D11.1+
    rom[300] = 11'b10011011001;	// +D12.1+
    rom[301] = 11'b11011001001;	// +D13.1+
    rom[302] = 11'b10111001001;	// +D14.1+
    rom[303] = 11'b01010001001;	// +D15.1-
    rom[304] = 11'b01001001001;	// +D16.1-
    rom[305] = 11'b11000111001;	// +D17.1+
    rom[306] = 11'b10100111001;	// +D18.1+
    rom[307] = 11'b11100101001;	// +D19.1+
    rom[308] = 11'b10010111001;	// +D20.1+
    rom[309] = 11'b11010101001;	// +D21.1+
    rom[310] = 11'b10110101001;	// +D22.1+
    rom[311] = 11'b00001011001;	// +D23.1-
    rom[312] = 11'b00011001001;	// +D24.1-
    rom[313] = 11'b11001101001;	// +D25.1+
    rom[314] = 11'b10101101001;	// +D26.1+
    rom[315] = 11'b00010011001;	// +D27.1-
    rom[316] = 11'b10011101001;	// +D28.1+
    rom[317] = 11'b00100011001;	// +D29.1-
    rom[318] = 11'b01000011001;	// +D30.1-
    rom[319] = 11'b00101001001;	// +D31.1-
    rom[320] = 11'b00110000101;	// +D00.2-
    rom[321] = 11'b01000100101;	// +D01.2-
    rom[322] = 11'b00100100101;	// +D02.2-
    rom[323] = 11'b11100010101;	// +D03.2+
    rom[324] = 11'b00010100101;	// +D04.2-
    rom[325] = 11'b11010010101;	// +D05.2+
    rom[326] = 11'b10110010101;	// +D06.2+
    rom[327] = 11'b10001110101;	// +D07.2+
    rom[328] = 11'b00001100101;	// +D08.2-
    rom[329] = 11'b11001010101;	// +D09.2+
    rom[330] = 11'b10101010101;	// +D10.2+
    rom[331] = 11'b11101000101;	// +D11.2+
    rom[332] = 11'b10011010101;	// +D12.2+
    rom[333] = 11'b11011000101;	// +D13.2+
    rom[334] = 11'b10111000101;	// +D14.2+
    rom[335] = 11'b01010000101;	// +D15.2-
    rom[336] = 11'b01001000101;	// +D16.2-
    rom[337] = 11'b11000110101;	// +D17.2+
    rom[338] = 11'b10100110101;	// +D18.2+
    rom[339] = 11'b11100100101;	// +D19.2+
    rom[340] = 11'b10010110101;	// +D20.2+
    rom[341] = 11'b11010100101;	// +D21.2+
    rom[342] = 11'b10110100101;	// +D22.2+
    rom[343] = 11'b00001010101;	// +D23.2-
    rom[344] = 11'b00011000101;	// +D24.2-
    rom[345] = 11'b11001100101;	// +D25.2+
    rom[346] = 11'b10101100101;	// +D26.2+
    rom[347] = 11'b00010010101;	// +D27.2-
    rom[348] = 11'b10011100101;	// +D28.2+
    rom[349] = 11'b00100010101;	// +D29.2-
    rom[350] = 11'b01000010101;	// +D30.2-
    rom[351] = 11'b00101000101;	// +D31.2-
    rom[352] = 11'b00110001100;	// +D00.3-
    rom[353] = 11'b01000101100;	// +D01.3-
    rom[354] = 11'b00100101100;	// +D02.3-
    rom[355] = 11'b11100010011;	// +D03.3+
    rom[356] = 11'b00010101100;	// +D04.3-
    rom[357] = 11'b11010010011;	// +D05.3+
    rom[358] = 11'b10110010011;	// +D06.3+
    rom[359] = 11'b10001110011;	// +D07.3+
    rom[360] = 11'b00001101100;	// +D08.3-
    rom[361] = 11'b11001010011;	// +D09.3+
    rom[362] = 11'b10101010011;	// +D10.3+
    rom[363] = 11'b11101000011;	// +D11.3+
    rom[364] = 11'b10011010011;	// +D12.3+
    rom[365] = 11'b11011000011;	// +D13.3+
    rom[366] = 11'b10111000011;	// +D14.3+
    rom[367] = 11'b01010001100;	// +D15.3-
    rom[368] = 11'b01001001100;	// +D16.3-
    rom[369] = 11'b11000110011;	// +D17.3+
    rom[370] = 11'b10100110011;	// +D18.3+
    rom[371] = 11'b11100100011;	// +D19.3+
    rom[372] = 11'b10010110011;	// +D20.3+
    rom[373] = 11'b11010100011;	// +D21.3+
    rom[374] = 11'b10110100011;	// +D22.3+
    rom[375] = 11'b00001011100;	// +D23.3-
    rom[376] = 11'b00011001100;	// +D24.3-
    rom[377] = 11'b11001100011;	// +D25.3+
    rom[378] = 11'b10101100011;	// +D26.3+
    rom[379] = 11'b00010011100;	// +D27.3-
    rom[380] = 11'b10011100011;	// +D28.3+
    rom[381] = 11'b00100011100;	// +D29.3-
    rom[382] = 11'b01000011100;	// +D30.3-
    rom[383] = 11'b00101001100;	// +D31.3-
    rom[384] = 11'b10110001101;	// +D00.4+
    rom[385] = 11'b11000101101;	// +D01.4+
    rom[386] = 11'b10100101101;	// +D02.4+
    rom[387] = 11'b01100010010;	// +D03.4-
    rom[388] = 11'b10010101101;	// +D04.4+
    rom[389] = 11'b01010010010;	// +D05.4-
    rom[390] = 11'b00110010010;	// +D06.4-
    rom[391] = 11'b00001110010;	// +D07.4-
    rom[392] = 11'b10001101101;	// +D08.4+
    rom[393] = 11'b01001010010;	// +D09.4-
    rom[394] = 11'b00101010010;	// +D10.4-
    rom[395] = 11'b01101000010;	// +D11.4-
    rom[396] = 11'b00011010010;	// +D12.4-
    rom[397] = 11'b01011000010;	// +D13.4-
    rom[398] = 11'b00111000010;	// +D14.4-
    rom[399] = 11'b11010001101;	// +D15.4+
    rom[400] = 11'b11001001101;	// +D16.4+
    rom[401] = 11'b01000110010;	// +D17.4-
    rom[402] = 11'b00100110010;	// +D18.4-
    rom[403] = 11'b01100100010;	// +D19.4-
    rom[404] = 11'b00010110010;	// +D20.4-
    rom[405] = 11'b01010100010;	// +D21.4-
    rom[406] = 11'b00110100010;	// +D22.4-
    rom[407] = 11'b10001011101;	// +D23.4+
    rom[408] = 11'b10011001101;	// +D24.4+
    rom[409] = 11'b01001100010;	// +D25.4-
    rom[410] = 11'b00101100010;	// +D26.4-
    rom[411] = 11'b10010011101;	// +D27.4+
    rom[412] = 11'b00011100010;	// +D28.4-
    rom[413] = 11'b10100011101;	// +D29.4+
    rom[414] = 11'b11000011101;	// +D30.4+
    rom[415] = 11'b10101001101;	// +D31.4+
    rom[416] = 11'b00110001010;	// +D00.5-
    rom[417] = 11'b01000101010;	// +D01.5-
    rom[418] = 11'b00100101010;	// +D02.5-
    rom[419] = 11'b11100011010;	// +D03.5+
    rom[420] = 11'b00010101010;	// +D04.5-
    rom[421] = 11'b11010011010;	// +D05.5+
    rom[422] = 11'b10110011010;	// +D06.5+
    rom[423] = 11'b10001111010;	// +D07.5+
    rom[424] = 11'b00001101010;	// +D08.5-
    rom[425] = 11'b11001011010;	// +D09.5+
    rom[426] = 11'b10101011010;	// +D10.5+
    rom[427] = 11'b11101001010;	// +D11.5+
    rom[428] = 11'b10011011010;	// +D12.5+
    rom[429] = 11'b11011001010;	// +D13.5+
    rom[430] = 11'b10111001010;	// +D14.5+
    rom[431] = 11'b01010001010;	// +D15.5-
    rom[432] = 11'b01001001010;	// +D16.5-
    rom[433] = 11'b11000111010;	// +D17.5+
    rom[434] = 11'b10100111010;	// +D18.5+
    rom[435] = 11'b11100101010;	// +D19.5+
    rom[436] = 11'b10010111010;	// +D20.5+
    rom[437] = 11'b11010101010;	// +D21.5+
    rom[438] = 11'b10110101010;	// +D22.5+
    rom[439] = 11'b00001011010;	// +D23.5-
    rom[440] = 11'b00011001010;	// +D24.5-
    rom[441] = 11'b11001101010;	// +D25.5+
    rom[442] = 11'b10101101010;	// +D26.5+
    rom[443] = 11'b00010011010;	// +D27.5-
    rom[444] = 11'b10011101010;	// +D28.5+
    rom[445] = 11'b00100011010;	// +D29.5-
    rom[446] = 11'b01000011010;	// +D30.5-
    rom[447] = 11'b00101001010;	// +D31.5-
    rom[448] = 11'b00110000110;	// +D00.6-
    rom[449] = 11'b01000100110;	// +D01.6-
    rom[450] = 11'b00100100110;	// +D02.6-
    rom[451] = 11'b11100010110;	// +D03.6+
    rom[452] = 11'b00010100110;	// +D04.6-
    rom[453] = 11'b11010010110;	// +D05.6+
    rom[454] = 11'b10110010110;	// +D06.6+
    rom[455] = 11'b10001110110;	// +D07.6+
    rom[456] = 11'b00001100110;	// +D08.6-
    rom[457] = 11'b11001010110;	// +D09.6+
    rom[458] = 11'b10101010110;	// +D10.6+
    rom[459] = 11'b11101000110;	// +D11.6+
    rom[460] = 11'b10011010110;	// +D12.6+
    rom[461] = 11'b11011000110;	// +D13.6+
    rom[462] = 11'b10111000110;	// +D14.6+
    rom[463] = 11'b01010000110;	// +D15.6-
    rom[464] = 11'b01001000110;	// +D16.6-
    rom[465] = 11'b11000110110;	// +D17.6+
    rom[466] = 11'b10100110110;	// +D18.6+
    rom[467] = 11'b11100100110;	// +D19.6+
    rom[468] = 11'b10010110110;	// +D20.6+
    rom[469] = 11'b11010100110;	// +D21.6+
    rom[470] = 11'b10110100110;	// +D22.6+
    rom[471] = 11'b00001010110;	// +D23.6-
    rom[472] = 11'b00011000110;	// +D24.6-
    rom[473] = 11'b11001100110;	// +D25.6+
    rom[474] = 11'b10101100110;	// +D26.6+
    rom[475] = 11'b00010010110;	// +D27.6-
    rom[476] = 11'b10011100110;	// +D28.6+
    rom[477] = 11'b00100010110;	// +D29.6-
    rom[478] = 11'b01000010110;	// +D30.6-
    rom[479] = 11'b00101000110;	// +D31.6-
    rom[480] = 11'b10110001110;	// +D00.7+
    rom[481] = 11'b11000101110;	// +D01.7+
    rom[482] = 11'b10100101110;	// +D02.7+
    rom[483] = 11'b01100010001;	// +D03.7-
    rom[484] = 11'b10010101110;	// +D04.7+
    rom[485] = 11'b01010010001;	// +D05.7-
    rom[486] = 11'b00110010001;	// +D06.7-
    rom[487] = 11'b00001110001;	// +D07.7-
    rom[488] = 11'b10001101110;	// +D08.7+
    rom[489] = 11'b01001010001;	// +D09.7-
    rom[490] = 11'b00101010001;	// +D10.7-
    rom[491] = 11'b01101001000;	// +D11.7-
    rom[492] = 11'b00011010001;	// +D12.7-
    rom[493] = 11'b01011001000;	// +D13.7-
    rom[494] = 11'b00111001000;	// +D14.7-
    rom[495] = 11'b11010001110;	// +D15.7+
    rom[496] = 11'b11001001110;	// +D16.7+
    rom[497] = 11'b01000110001;	// +D17.7-
    rom[498] = 11'b00100110001;	// +D18.7-
    rom[499] = 11'b01100100001;	// +D19.7-
    rom[500] = 11'b00010110001;	// +D20.7-
    rom[501] = 11'b01010100001;	// +D21.7-
    rom[502] = 11'b00110100001;	// +D22.7-
    rom[503] = 11'b10001011110;	// +D23.7+
    rom[504] = 11'b10011001110;	// +D24.7+
    rom[505] = 11'b01001100001;	// +D25.7-
    rom[506] = 11'b00101100001;	// +D26.7-
    rom[507] = 11'b10010011110;	// +D27.7+
    rom[508] = 11'b00011100001;	// +D28.7-
    rom[509] = 11'b10100011110;	// +D29.7+
    rom[510] = 11'b11000011110;	// +D30.7+
    rom[511] = 11'b10101001110;	// +D31.7+
    rom[512] = 11'b01001110100;	// -K00.0-
    rom[513] = 11'b00111010100;	// -K01.0-
    rom[514] = 11'b01011010100;	// -K02.0-
    rom[515] = 11'b11100011011;	// -K03.0+
    rom[516] = 11'b01101010100;	// -K04.0-
    rom[517] = 11'b11010011011;	// -K05.0+
    rom[518] = 11'b10110011011;	// -K06.0+
    rom[519] = 11'b11110001011;	// -K07.0+
    rom[520] = 11'b01110010100;	// -K08.0-
    rom[521] = 11'b11001011011;	// -K09.0+
    rom[522] = 11'b10101011011;	// -K10.0+
    rom[523] = 11'b11101001011;	// -K11.0+
    rom[524] = 11'b10011011011;	// -K12.0+
    rom[525] = 11'b11011001011;	// -K13.0+
    rom[526] = 11'b10111001011;	// -K14.0+
    rom[527] = 11'b00101110100;	// -K15.0-
    rom[528] = 11'b00110110100;	// -K16.0-
    rom[529] = 11'b11000111011;	// -K17.0+
    rom[530] = 11'b10100111011;	// -K18.0+
    rom[531] = 11'b11100101011;	// -K19.0+
    rom[532] = 11'b10010111011;	// -K20.0+
    rom[533] = 11'b11010101011;	// -K21.0+
    rom[534] = 11'b10110101011;	// -K22.0+
    rom[535] = 11'b01110100100;	// -K23.0-
    rom[536] = 11'b01100110100;	// -K24.0-
    rom[537] = 11'b11001101011;	// -K25.0+
    rom[538] = 11'b10101101011;	// -K26.0+
    rom[539] = 11'b01101100100;	// -K27.0-
    rom[540] = 11'b00011110100;	// -K28.0-
    rom[541] = 11'b01011100100;	// -K29.0-
    rom[542] = 11'b00111100100;	// -K30.0-
    rom[543] = 11'b01010110100;	// -K31.0-
    rom[544] = 11'b11001111001;	// -K00.1+
    rom[545] = 11'b10111011001;	// -K01.1+
    rom[546] = 11'b11011011001;	// -K02.1+
    rom[547] = 11'b01100010110;	// -K03.1-
    rom[548] = 11'b11101011001;	// -K04.1+
    rom[549] = 11'b01010010110;	// -K05.1-
    rom[550] = 11'b00110010110;	// -K06.1-
    rom[551] = 11'b01110000110;	// -K07.1-
    rom[552] = 11'b11110011001;	// -K08.1+
    rom[553] = 11'b01001010110;	// -K09.1-
    rom[554] = 11'b00101010110;	// -K10.1-
    rom[555] = 11'b01101000110;	// -K11.1-
    rom[556] = 11'b00011010110;	// -K12.1-
    rom[557] = 11'b01011000110;	// -K13.1-
    rom[558] = 11'b00111000110;	// -K14.1-
    rom[559] = 11'b10101111001;	// -K15.1+
    rom[560] = 11'b10110111001;	// -K16.1+
    rom[561] = 11'b01000110110;	// -K17.1-
    rom[562] = 11'b00100110110;	// -K18.1-
    rom[563] = 11'b01100100110;	// -K19.1-
    rom[564] = 11'b00010110110;	// -K20.1-
    rom[565] = 11'b01010100110;	// -K21.1-
    rom[566] = 11'b00110100110;	// -K22.1-
    rom[567] = 11'b11110101001;	// -K23.1+
    rom[568] = 11'b11100111001;	// -K24.1+
    rom[569] = 11'b01001100110;	// -K25.1-
    rom[570] = 11'b00101100110;	// -K26.1-
    rom[571] = 11'b11101101001;	// -K27.1+
    rom[572] = 11'b10011111001;	// -K28.1+
    rom[573] = 11'b11011101001;	// -K29.1+
    rom[574] = 11'b10111101001;	// -K30.1+
    rom[575] = 11'b11010111001;	// -K31.1+
    rom[576] = 11'b11001110101;	// -K00.2+
    rom[577] = 11'b10111010101;	// -K01.2+
    rom[578] = 11'b11011010101;	// -K02.2+
    rom[579] = 11'b01100011010;	// -K03.2-
    rom[580] = 11'b11101010101;	// -K04.2+
    rom[581] = 11'b01010011010;	// -K05.2-
    rom[582] = 11'b00110011010;	// -K06.2-
    rom[583] = 11'b01110001010;	// -K07.2-
    rom[584] = 11'b11110010101;	// -K08.2+
    rom[585] = 11'b01001011010;	// -K09.2-
    rom[586] = 11'b00101011010;	// -K10.2-
    rom[587] = 11'b01101001010;	// -K11.2-
    rom[588] = 11'b00011011010;	// -K12.2-
    rom[589] = 11'b01011001010;	// -K13.2-
    rom[590] = 11'b00111001010;	// -K14.2-
    rom[591] = 11'b10101110101;	// -K15.2+
    rom[592] = 11'b10110110101;	// -K16.2+
    rom[593] = 11'b01000111010;	// -K17.2-
    rom[594] = 11'b00100111010;	// -K18.2-
    rom[595] = 11'b01100101010;	// -K19.2-
    rom[596] = 11'b00010111010;	// -K20.2-
    rom[597] = 11'b01010101010;	// -K21.2-
    rom[598] = 11'b00110101010;	// -K22.2-
    rom[599] = 11'b11110100101;	// -K23.2+
    rom[600] = 11'b11100110101;	// -K24.2+
    rom[601] = 11'b01001101010;	// -K25.2-
    rom[602] = 11'b00101101010;	// -K26.2-
    rom[603] = 11'b11101100101;	// -K27.2+
    rom[604] = 11'b10011110101;	// -K28.2+
    rom[605] = 11'b11011100101;	// -K29.2+
    rom[606] = 11'b10111100101;	// -K30.2+
    rom[607] = 11'b11010110101;	// -K31.2+
    rom[608] = 11'b11001110011;	// -K00.3+
    rom[609] = 11'b10111010011;	// -K01.3+
    rom[610] = 11'b11011010011;	// -K02.3+
    rom[611] = 11'b01100011100;	// -K03.3-
    rom[612] = 11'b11101010011;	// -K04.3+
    rom[613] = 11'b01010011100;	// -K05.3-
    rom[614] = 11'b00110011100;	// -K06.3-
    rom[615] = 11'b01110001100;	// -K07.3-
    rom[616] = 11'b11110010011;	// -K08.3+
    rom[617] = 11'b01001011100;	// -K09.3-
    rom[618] = 11'b00101011100;	// -K10.3-
    rom[619] = 11'b01101001100;	// -K11.3-
    rom[620] = 11'b00011011100;	// -K12.3-
    rom[621] = 11'b01011001100;	// -K13.3-
    rom[622] = 11'b00111001100;	// -K14.3-
    rom[623] = 11'b10101110011;	// -K15.3+
    rom[624] = 11'b10110110011;	// -K16.3+
    rom[625] = 11'b01000111100;	// -K17.3-
    rom[626] = 11'b00100111100;	// -K18.3-
    rom[627] = 11'b01100101100;	// -K19.3-
    rom[628] = 11'b00010111100;	// -K20.3-
    rom[629] = 11'b01010101100;	// -K21.3-
    rom[630] = 11'b00110101100;	// -K22.3-
    rom[631] = 11'b11110100011;	// -K23.3+
    rom[632] = 11'b11100110011;	// -K24.3+
    rom[633] = 11'b01001101100;	// -K25.3-
    rom[634] = 11'b00101101100;	// -K26.3-
    rom[635] = 11'b11101100011;	// -K27.3+
    rom[636] = 11'b10011110011;	// -K28.3+
    rom[637] = 11'b11011100011;	// -K29.3+
    rom[638] = 11'b10111100011;	// -K30.3+
    rom[639] = 11'b11010110011;	// -K31.3+
    rom[640] = 11'b01001110010;	// -K00.4-
    rom[641] = 11'b00111010010;	// -K01.4-
    rom[642] = 11'b01011010010;	// -K02.4-
    rom[643] = 11'b11100011101;	// -K03.4+
    rom[644] = 11'b01101010010;	// -K04.4-
    rom[645] = 11'b11010011101;	// -K05.4+
    rom[646] = 11'b10110011101;	// -K06.4+
    rom[647] = 11'b11110001101;	// -K07.4+
    rom[648] = 11'b01110010010;	// -K08.4-
    rom[649] = 11'b11001011101;	// -K09.4+
    rom[650] = 11'b10101011101;	// -K10.4+
    rom[651] = 11'b11101001101;	// -K11.4+
    rom[652] = 11'b10011011101;	// -K12.4+
    rom[653] = 11'b11011001101;	// -K13.4+
    rom[654] = 11'b10111001101;	// -K14.4+
    rom[655] = 11'b00101110010;	// -K15.4-
    rom[656] = 11'b00110110010;	// -K16.4-
    rom[657] = 11'b11000111101;	// -K17.4+
    rom[658] = 11'b10100111101;	// -K18.4+
    rom[659] = 11'b11100101101;	// -K19.4+
    rom[660] = 11'b10010111101;	// -K20.4+
    rom[661] = 11'b11010101101;	// -K21.4+
    rom[662] = 11'b10110101101;	// -K22.4+
    rom[663] = 11'b01110100010;	// -K23.4-
    rom[664] = 11'b01100110010;	// -K24.4-
    rom[665] = 11'b11001101101;	// -K25.4+
    rom[666] = 11'b10101101101;	// -K26.4+
    rom[667] = 11'b01101100010;	// -K27.4-
    rom[668] = 11'b00011110010;	// -K28.4-
    rom[669] = 11'b01011100010;	// -K29.4-
    rom[670] = 11'b00111100010;	// -K30.4-
    rom[671] = 11'b01010110010;	// -K31.4-
    rom[672] = 11'b11001111010;	// -K00.5+
    rom[673] = 11'b10111011010;	// -K01.5+
    rom[674] = 11'b11011011010;	// -K02.5+
    rom[675] = 11'b01100010101;	// -K03.5-
    rom[676] = 11'b11101011010;	// -K04.5+
    rom[677] = 11'b01010010101;	// -K05.5-
    rom[678] = 11'b00110010101;	// -K06.5-
    rom[679] = 11'b01110000101;	// -K07.5-
    rom[680] = 11'b11110011010;	// -K08.5+
    rom[681] = 11'b01001010101;	// -K09.5-
    rom[682] = 11'b00101010101;	// -K10.5-
    rom[683] = 11'b01101000101;	// -K11.5-
    rom[684] = 11'b00011010101;	// -K12.5-
    rom[685] = 11'b01011000101;	// -K13.5-
    rom[686] = 11'b00111000101;	// -K14.5-
    rom[687] = 11'b10101111010;	// -K15.5+
    rom[688] = 11'b10110111010;	// -K16.5+
    rom[689] = 11'b01000110101;	// -K17.5-
    rom[690] = 11'b00100110101;	// -K18.5-
    rom[691] = 11'b01100100101;	// -K19.5-
    rom[692] = 11'b00010110101;	// -K20.5-
    rom[693] = 11'b01010100101;	// -K21.5-
    rom[694] = 11'b00110100101;	// -K22.5-
    rom[695] = 11'b11110101010;	// -K23.5+
    rom[696] = 11'b11100111010;	// -K24.5+
    rom[697] = 11'b01001100101;	// -K25.5-
    rom[698] = 11'b00101100101;	// -K26.5-
    rom[699] = 11'b11101101010;	// -K27.5+
    rom[700] = 11'b10011111010;	// -K28.5+
    rom[701] = 11'b11011101010;	// -K29.5+
    rom[702] = 11'b10111101010;	// -K30.5+
    rom[703] = 11'b11010111010;	// -K31.5+
    rom[704] = 11'b11001110110;	// -K00.6+
    rom[705] = 11'b10111010110;	// -K01.6+
    rom[706] = 11'b11011010110;	// -K02.6+
    rom[707] = 11'b01100011001;	// -K03.6-
    rom[708] = 11'b11101010110;	// -K04.6+
    rom[709] = 11'b01010011001;	// -K05.6-
    rom[710] = 11'b00110011001;	// -K06.6-
    rom[711] = 11'b01110001001;	// -K07.6-
    rom[712] = 11'b11110010110;	// -K08.6+
    rom[713] = 11'b01001011001;	// -K09.6-
    rom[714] = 11'b00101011001;	// -K10.6-
    rom[715] = 11'b01101001001;	// -K11.6-
    rom[716] = 11'b00011011001;	// -K12.6-
    rom[717] = 11'b01011001001;	// -K13.6-
    rom[718] = 11'b00111001001;	// -K14.6-
    rom[719] = 11'b10101110110;	// -K15.6+
    rom[720] = 11'b10110110110;	// -K16.6+
    rom[721] = 11'b01000111001;	// -K17.6-
    rom[722] = 11'b00100111001;	// -K18.6-
    rom[723] = 11'b01100101001;	// -K19.6-
    rom[724] = 11'b00010111001;	// -K20.6-
    rom[725] = 11'b01010101001;	// -K21.6-
    rom[726] = 11'b00110101001;	// -K22.6-
    rom[727] = 11'b11110100110;	// -K23.6+
    rom[728] = 11'b11100110110;	// -K24.6+
    rom[729] = 11'b01001101001;	// -K25.6-
    rom[730] = 11'b00101101001;	// -K26.6-
    rom[731] = 11'b11101100110;	// -K27.6+
    rom[732] = 11'b10011110110;	// -K28.6+
    rom[733] = 11'b11011100110;	// -K29.6+
    rom[734] = 11'b10111100110;	// -K30.6+
    rom[735] = 11'b11010110110;	// -K31.6+
    rom[736] = 11'b01001111000;	// -K00.7-
    rom[737] = 11'b00111011000;	// -K01.7-
    rom[738] = 11'b01011011000;	// -K02.7-
    rom[739] = 11'b11100010111;	// -K03.7+
    rom[740] = 11'b01101011000;	// -K04.7-
    rom[741] = 11'b11010010111;	// -K05.7+
    rom[742] = 11'b10110010111;	// -K06.7+
    rom[743] = 11'b11110000111;	// -K07.7+
    rom[744] = 11'b01110011000;	// -K08.7-
    rom[745] = 11'b11001010111;	// -K09.7+
    rom[746] = 11'b10101010111;	// -K10.7+
    rom[747] = 11'b11101000111;	// -K11.7+
    rom[748] = 11'b10011010111;	// -K12.7+
    rom[749] = 11'b11011000111;	// -K13.7+
    rom[750] = 11'b10111000111;	// -K14.7+
    rom[751] = 11'b00101111000;	// -K15.7-
    rom[752] = 11'b00110111000;	// -K16.7-
    rom[753] = 11'b11000110111;	// -K17.7+
    rom[754] = 11'b10100110111;	// -K18.7+
    rom[755] = 11'b11100100111;	// -K19.7+
    rom[756] = 11'b10010110111;	// -K20.7+
    rom[757] = 11'b11010100111;	// -K21.7+
    rom[758] = 11'b10110100111;	// -K22.7+
    rom[759] = 11'b01110101000;	// -K23.7-
    rom[760] = 11'b01100111000;	// -K24.7-
    rom[761] = 11'b11001100111;	// -K25.7+
    rom[762] = 11'b10101100111;	// -K26.7+
    rom[763] = 11'b01101101000;	// -K27.7-
    rom[764] = 11'b00011111000;	// -K28.7-
    rom[765] = 11'b01011101000;	// -K29.7-
    rom[766] = 11'b00111101000;	// -K30.7-
    rom[767] = 11'b01010111000;	// -K31.7-
    rom[768] = 11'b10110001011;	// +K00.0+
    rom[769] = 11'b11000101011;	// +K01.0+
    rom[770] = 11'b10100101011;	// +K02.0+
    rom[771] = 11'b01100010100;	// +K03.0-
    rom[772] = 11'b10010101011;	// +K04.0+
    rom[773] = 11'b01010010100;	// +K05.0-
    rom[774] = 11'b00110010100;	// +K06.0-
    rom[775] = 11'b00001110100;	// +K07.0-
    rom[776] = 11'b10001101011;	// +K08.0+
    rom[777] = 11'b01001010100;	// +K09.0-
    rom[778] = 11'b00101010100;	// +K10.0-
    rom[779] = 11'b01101000100;	// +K11.0-
    rom[780] = 11'b00011010100;	// +K12.0-
    rom[781] = 11'b01011000100;	// +K13.0-
    rom[782] = 11'b00111000100;	// +K14.0-
    rom[783] = 11'b11010001011;	// +K15.0+
    rom[784] = 11'b11001001011;	// +K16.0+
    rom[785] = 11'b01000110100;	// +K17.0-
    rom[786] = 11'b00100110100;	// +K18.0-
    rom[787] = 11'b01100100100;	// +K19.0-
    rom[788] = 11'b00010110100;	// +K20.0-
    rom[789] = 11'b01010100100;	// +K21.0-
    rom[790] = 11'b00110100100;	// +K22.0-
    rom[791] = 11'b10001011011;	// +K23.0+
    rom[792] = 11'b10011001011;	// +K24.0+
    rom[793] = 11'b01001100100;	// +K25.0-
    rom[794] = 11'b00101100100;	// +K26.0-
    rom[795] = 11'b10010011011;	// +K27.0+
    rom[796] = 11'b11100001011;	// +K28.0+
    rom[797] = 11'b10100011011;	// +K29.0+
    rom[798] = 11'b11000011011;	// +K30.0+
    rom[799] = 11'b10101001011;	// +K31.0+
    rom[800] = 11'b00110000110;	// +K00.1-
    rom[801] = 11'b01000100110;	// +K01.1-
    rom[802] = 11'b00100100110;	// +K02.1-
    rom[803] = 11'b11100011001;	// +K03.1+
    rom[804] = 11'b00010100110;	// +K04.1-
    rom[805] = 11'b11010011001;	// +K05.1+
    rom[806] = 11'b10110011001;	// +K06.1+
    rom[807] = 11'b10001111001;	// +K07.1+
    rom[808] = 11'b00001100110;	// +K08.1-
    rom[809] = 11'b11001011001;	// +K09.1+
    rom[810] = 11'b10101011001;	// +K10.1+
    rom[811] = 11'b11101001001;	// +K11.1+
    rom[812] = 11'b10011011001;	// +K12.1+
    rom[813] = 11'b11011001001;	// +K13.1+
    rom[814] = 11'b10111001001;	// +K14.1+
    rom[815] = 11'b01010000110;	// +K15.1-
    rom[816] = 11'b01001000110;	// +K16.1-
    rom[817] = 11'b11000111001;	// +K17.1+
    rom[818] = 11'b10100111001;	// +K18.1+
    rom[819] = 11'b11100101001;	// +K19.1+
    rom[820] = 11'b10010111001;	// +K20.1+
    rom[821] = 11'b11010101001;	// +K21.1+
    rom[822] = 11'b10110101001;	// +K22.1+
    rom[823] = 11'b00001010110;	// +K23.1-
    rom[824] = 11'b00011000110;	// +K24.1-
    rom[825] = 11'b11001101001;	// +K25.1+
    rom[826] = 11'b10101101001;	// +K26.1+
    rom[827] = 11'b00010010110;	// +K27.1-
    rom[828] = 11'b01100000110;	// +K28.1-
    rom[829] = 11'b00100010110;	// +K29.1-
    rom[830] = 11'b01000010110;	// +K30.1-
    rom[831] = 11'b00101000110;	// +K31.1-
    rom[832] = 11'b00110001010;	// +K00.2-
    rom[833] = 11'b01000101010;	// +K01.2-
    rom[834] = 11'b00100101010;	// +K02.2-
    rom[835] = 11'b11100010101;	// +K03.2+
    rom[836] = 11'b00010101010;	// +K04.2-
    rom[837] = 11'b11010010101;	// +K05.2+
    rom[838] = 11'b10110010101;	// +K06.2+
    rom[839] = 11'b10001110101;	// +K07.2+
    rom[840] = 11'b00001101010;	// +K08.2-
    rom[841] = 11'b11001010101;	// +K09.2+
    rom[842] = 11'b10101010101;	// +K10.2+
    rom[843] = 11'b11101000101;	// +K11.2+
    rom[844] = 11'b10011010101;	// +K12.2+
    rom[845] = 11'b11011000101;	// +K13.2+
    rom[846] = 11'b10111000101;	// +K14.2+
    rom[847] = 11'b01010001010;	// +K15.2-
    rom[848] = 11'b01001001010;	// +K16.2-
    rom[849] = 11'b11000110101;	// +K17.2+
    rom[850] = 11'b10100110101;	// +K18.2+
    rom[851] = 11'b11100100101;	// +K19.2+
    rom[852] = 11'b10010110101;	// +K20.2+
    rom[853] = 11'b11010100101;	// +K21.2+
    rom[854] = 11'b10110100101;	// +K22.2+
    rom[855] = 11'b00001011010;	// +K23.2-
    rom[856] = 11'b00011001010;	// +K24.2-
    rom[857] = 11'b11001100101;	// +K25.2+
    rom[858] = 11'b10101100101;	// +K26.2+
    rom[859] = 11'b00010011010;	// +K27.2-
    rom[860] = 11'b01100001010;	// +K28.2-
    rom[861] = 11'b00100011010;	// +K29.2-
    rom[862] = 11'b01000011010;	// +K30.2-
    rom[863] = 11'b00101001010;	// +K31.2-
    rom[864] = 11'b00110001100;	// +K00.3-
    rom[865] = 11'b01000101100;	// +K01.3-
    rom[866] = 11'b00100101100;	// +K02.3-
    rom[867] = 11'b11100010011;	// +K03.3+
    rom[868] = 11'b00010101100;	// +K04.3-
    rom[869] = 11'b11010010011;	// +K05.3+
    rom[870] = 11'b10110010011;	// +K06.3+
    rom[871] = 11'b10001110011;	// +K07.3+
    rom[872] = 11'b00001101100;	// +K08.3-
    rom[873] = 11'b11001010011;	// +K09.3+
    rom[874] = 11'b10101010011;	// +K10.3+
    rom[875] = 11'b11101000011;	// +K11.3+
    rom[876] = 11'b10011010011;	// +K12.3+
    rom[877] = 11'b11011000011;	// +K13.3+
    rom[878] = 11'b10111000011;	// +K14.3+
    rom[879] = 11'b01010001100;	// +K15.3-
    rom[880] = 11'b01001001100;	// +K16.3-
    rom[881] = 11'b11000110011;	// +K17.3+
    rom[882] = 11'b10100110011;	// +K18.3+
    rom[883] = 11'b11100100011;	// +K19.3+
    rom[884] = 11'b10010110011;	// +K20.3+
    rom[885] = 11'b11010100011;	// +K21.3+
    rom[886] = 11'b10110100011;	// +K22.3+
    rom[887] = 11'b00001011100;	// +K23.3-
    rom[888] = 11'b00011001100;	// +K24.3-
    rom[889] = 11'b11001100011;	// +K25.3+
    rom[890] = 11'b10101100011;	// +K26.3+
    rom[891] = 11'b00010011100;	// +K27.3-
    rom[892] = 11'b01100001100;	// +K28.3-
    rom[893] = 11'b00100011100;	// +K29.3-
    rom[894] = 11'b01000011100;	// +K30.3-
    rom[895] = 11'b00101001100;	// +K31.3-
    rom[896] = 11'b10110001101;	// +K00.4+
    rom[897] = 11'b11000101101;	// +K01.4+
    rom[898] = 11'b10100101101;	// +K02.4+
    rom[899] = 11'b01100010010;	// +K03.4-
    rom[900] = 11'b10010101101;	// +K04.4+
    rom[901] = 11'b01010010010;	// +K05.4-
    rom[902] = 11'b00110010010;	// +K06.4-
    rom[903] = 11'b00001110010;	// +K07.4-
    rom[904] = 11'b10001101101;	// +K08.4+
    rom[905] = 11'b01001010010;	// +K09.4-
    rom[906] = 11'b00101010010;	// +K10.4-
    rom[907] = 11'b01101000010;	// +K11.4-
    rom[908] = 11'b00011010010;	// +K12.4-
    rom[909] = 11'b01011000010;	// +K13.4-
    rom[910] = 11'b00111000010;	// +K14.4-
    rom[911] = 11'b11010001101;	// +K15.4+
    rom[912] = 11'b11001001101;	// +K16.4+
    rom[913] = 11'b01000110010;	// +K17.4-
    rom[914] = 11'b00100110010;	// +K18.4-
    rom[915] = 11'b01100100010;	// +K19.4-
    rom[916] = 11'b00010110010;	// +K20.4-
    rom[917] = 11'b01010100010;	// +K21.4-
    rom[918] = 11'b00110100010;	// +K22.4-
    rom[919] = 11'b10001011101;	// +K23.4+
    rom[920] = 11'b10011001101;	// +K24.4+
    rom[921] = 11'b01001100010;	// +K25.4-
    rom[922] = 11'b00101100010;	// +K26.4-
    rom[923] = 11'b10010011101;	// +K27.4+
    rom[924] = 11'b11100001101;	// +K28.4+
    rom[925] = 11'b10100011101;	// +K29.4+
    rom[926] = 11'b11000011101;	// +K30.4+
    rom[927] = 11'b10101001101;	// +K31.4+
    rom[928] = 11'b00110000101;	// +K00.5-
    rom[929] = 11'b01000100101;	// +K01.5-
    rom[930] = 11'b00100100101;	// +K02.5-
    rom[931] = 11'b11100011010;	// +K03.5+
    rom[932] = 11'b00010100101;	// +K04.5-
    rom[933] = 11'b11010011010;	// +K05.5+
    rom[934] = 11'b10110011010;	// +K06.5+
    rom[935] = 11'b10001111010;	// +K07.5+
    rom[936] = 11'b00001100101;	// +K08.5-
    rom[937] = 11'b11001011010;	// +K09.5+
    rom[938] = 11'b10101011010;	// +K10.5+
    rom[939] = 11'b11101001010;	// +K11.5+
    rom[940] = 11'b10011011010;	// +K12.5+
    rom[941] = 11'b11011001010;	// +K13.5+
    rom[942] = 11'b10111001010;	// +K14.5+
    rom[943] = 11'b01010000101;	// +K15.5-
    rom[944] = 11'b01001000101;	// +K16.5-
    rom[945] = 11'b11000111010;	// +K17.5+
    rom[946] = 11'b10100111010;	// +K18.5+
    rom[947] = 11'b11100101010;	// +K19.5+
    rom[948] = 11'b10010111010;	// +K20.5+
    rom[949] = 11'b11010101010;	// +K21.5+
    rom[950] = 11'b10110101010;	// +K22.5+
    rom[951] = 11'b00001010101;	// +K23.5-
    rom[952] = 11'b00011000101;	// +K24.5-
    rom[953] = 11'b11001101010;	// +K25.5+
    rom[954] = 11'b10101101010;	// +K26.5+
    rom[955] = 11'b00010010101;	// +K27.5-
    rom[956] = 11'b01100000101;	// +K28.5-
    rom[957] = 11'b00100010101;	// +K29.5-
    rom[958] = 11'b01000010101;	// +K30.5-
    rom[959] = 11'b00101000101;	// +K31.5-
    rom[960] = 11'b00110001001;	// +K00.6-
    rom[961] = 11'b01000101001;	// +K01.6-
    rom[962] = 11'b00100101001;	// +K02.6-
    rom[963] = 11'b11100010110;	// +K03.6+
    rom[964] = 11'b00010101001;	// +K04.6-
    rom[965] = 11'b11010010110;	// +K05.6+
    rom[966] = 11'b10110010110;	// +K06.6+
    rom[967] = 11'b10001110110;	// +K07.6+
    rom[968] = 11'b00001101001;	// +K08.6-
    rom[969] = 11'b11001010110;	// +K09.6+
    rom[970] = 11'b10101010110;	// +K10.6+
    rom[971] = 11'b11101000110;	// +K11.6+
    rom[972] = 11'b10011010110;	// +K12.6+
    rom[973] = 11'b11011000110;	// +K13.6+
    rom[974] = 11'b10111000110;	// +K14.6+
    rom[975] = 11'b01010001001;	// +K15.6-
    rom[976] = 11'b01001001001;	// +K16.6-
    rom[977] = 11'b11000110110;	// +K17.6+
    rom[978] = 11'b10100110110;	// +K18.6+
    rom[979] = 11'b11100100110;	// +K19.6+
    rom[980] = 11'b10010110110;	// +K20.6+
    rom[981] = 11'b11010100110;	// +K21.6+
    rom[982] = 11'b10110100110;	// +K22.6+
    rom[983] = 11'b00001011001;	// +K23.6-
    rom[984] = 11'b00011001001;	// +K24.6-
    rom[985] = 11'b11001100110;	// +K25.6+
    rom[986] = 11'b10101100110;	// +K26.6+
    rom[987] = 11'b00010011001;	// +K27.6-
    rom[988] = 11'b01100001001;	// +K28.6-
    rom[989] = 11'b00100011001;	// +K29.6-
    rom[990] = 11'b01000011001;	// +K30.6-
    rom[991] = 11'b00101001001;	// +K31.6-
    rom[992] = 11'b10110000111;	// +K00.7+
    rom[993] = 11'b11000100111;	// +K01.7+
    rom[994] = 11'b10100100111;	// +K02.7+
    rom[995] = 11'b01100011000;	// +K03.7-
    rom[996] = 11'b10010100111;	// +K04.7+
    rom[997] = 11'b01010011000;	// +K05.7-
    rom[998] = 11'b00110011000;	// +K06.7-
    rom[999] = 11'b00001111000;	// +K07.7-
    rom[1000] = 11'b10001100111;	// +K08.7+
    rom[1001] = 11'b01001011000;	// +K09.7-
    rom[1002] = 11'b00101011000;	// +K10.7-
    rom[1003] = 11'b01101001000;	// +K11.7-
    rom[1004] = 11'b00011011000;	// +K12.7-
    rom[1005] = 11'b01011001000;	// +K13.7-
    rom[1006] = 11'b00111001000;	// +K14.7-
    rom[1007] = 11'b11010000111;	// +K15.7+
    rom[1008] = 11'b11001000111;	// +K16.7+
    rom[1009] = 11'b01000111000;	// +K17.7-
    rom[1010] = 11'b00100111000;	// +K18.7-
    rom[1011] = 11'b01100101000;	// +K19.7-
    rom[1012] = 11'b00010111000;	// +K20.7-
    rom[1013] = 11'b01010101000;	// +K21.7-
    rom[1014] = 11'b00110101000;	// +K22.7-
    rom[1015] = 11'b10001010111;	// +K23.7+
    rom[1016] = 11'b10011000111;	// +K24.7+
    rom[1017] = 11'b01001101000;	// +K25.7-
    rom[1018] = 11'b00101101000;	// +K26.7-
    rom[1019] = 11'b10010010111;	// +K27.7+
    rom[1020] = 11'b11100000111;	// +K28.7+
    rom[1021] = 11'b10100010111;	// +K29.7+
    rom[1022] = 11'b11000010111;	// +K30.7+
    rom[1023] = 11'b10101000111;	// +K31.7+
  end

endmodule : encoder_8b10b
